class test extends uvm_test;
  `uvm_component_utils(test)
  
  function new(input string inst = "TEST", uvm_component c);
    super.new(inst,c);
    endfunction
  
  sequence_random gen;
  env e;
  
  
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    gen=sequence_random::type_id::create("gen",this);
    e =env::type_id::create("e",this);
  endfunction
  
  virtual task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    gen.start(e.a.seqr);
    phase.drop_objection(this);
  endtask
endclass
